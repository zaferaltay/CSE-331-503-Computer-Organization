module shiftLeft2_32Bit(input1,output1);

input [31:0]input1;
output [31:0] output1;


assign output1[31]=input1[29];
assign output1[30]=input1[28];
assign output1[29]=input1[27];
assign output1[28]=input1[26];
assign output1[27]=input1[25];
assign output1[26]=input1[24];
assign output1[25]=input1[23];
assign output1[24]=input1[22];
assign output1[23]=input1[21];
assign output1[22]=input1[20];
assign output1[21]=input1[19];
assign output1[20]=input1[18];
assign output1[19]=input1[17];
assign output1[18]=input1[16];
assign output1[17]=input1[15];
assign output1[16]=input1[14];
assign output1[15]=input1[13];
assign output1[14]=input1[12];
assign output1[13]=input1[11];
assign output1[12]=input1[10];
assign output1[11]=input1[9];
assign output1[10]=input1[8];
assign output1[9]=input1[7];
assign output1[8]=input1[6];
assign output1[7]=input1[5];
assign output1[6]=input1[4];
assign output1[5]=input1[3];
assign output1[4]=input1[2];
assign output1[3]=input1[1];
assign output1[2]=input1[0];
assign output1[1]=1'b0;
assign output1[0]=1'b0;




endmodule